`timescale 1ns / 1ps

module inst_mem (
    input  logic [31:0] inst_read_addr,
    output logic [31:0] inst_code
);
    logic [31:0] rom[0:1023]; // byte align 256*4

    initial begin
        $readmemh("code.mem", rom);
        // for(int i = 0; i<64; i++) begin
        //     rom[i] = 32'hffff_0000+i;
        // end

        // rom[0] = 32'b0000000_00100_01000_000_00101_0110011;  // add x5, x8, x4    12
        // rom[1] = 32'b0100000_01001_01000_000_00111_0110011;  // sub x7, x8, x9    -1

        // // B-type
        // // 32'b imm(7bit) rs2(5bit) _ rs1(5bit) _ funct3(3bit) _ imm (5bit) _ opcode(7'b1100011)
        // rom[2] =  32'b0000000_00010_00010_000_01000_1100011; // BEQ x2, x2, 8
        // rom[4] =  32'b0000000_00010_00001_001_01000_1100011; // BNE x1, x2, 8
        // rom[6] =  32'b0000000_00010_00001_100_01000_1100011; // BLT x1, x2, 8 (signed) 
        // rom[8] =  32'b0000000_00001_00010_101_01000_1100011; // BGE x2, x1, 8 (signed)     0
        // rom[10] = 32'b0000000_00010_00001_110_01000_1100011; // BLTU x1, x2, 8 (unsigned  1
        // rom[12] = 32'b0000000_00001_00010_111_01000_1100011; // BGEU x2, x1, 8 (unsigned)  0

        // // S-type
        // // 32'b imm(7bit) _ rs2(5bit) _ rs1(5bit) _ funct3(3bit) _ imm (5bit) opcode(7'b0100011)
        // rom[13] = 32'b0000000_01000_00000_000_00000_0100011;  // sb x2, 0(x0)
        // rom[14] = 32'b0000000_00100_00000_001_00010_0100011;  // sh x2, 2(x0)
        // rom[15] = 32'b0000000_00010_00000_010_00100_0100011;  // sw x2, 4(x0)

        // // I-type LOAD
        // rom[16] = 32'b000000000100_00001_000_00101_0000011;  // LB  x5, 4(x1)
        // rom[17] = 32'b000000001000_00001_001_00101_0000011;  // LH  x5, 8(x1)
        // rom[18] = 32'b000000001100_00001_010_00101_0000011;  // LW  x5, 12(x1)
        // rom[19] = 32'b000000010000_00001_100_00101_0000011;  // LBU x5, 16(x1)
        // rom[20] = 32'b000000010100_00001_101_00101_0000011;  // LHU x5, 20(x1)

        // // I-type ALU Immediate
        // rom[21] = 32'h00C30413;  // addi x8, x6, 12
        // rom[22] = 32'b000000000101_00110_010_01001_0010011;  // slti x9, x6, 5
        // rom[23] = 32'b000000000111_00110_111_01010_0010011;  // andi x10, x6, 7
        // rom[24] = 32'b000000001010_00110_110_01011_0010011;  // ori  x11, x6, 10
        // rom[25] = 32'b000000001100_00110_100_01100_0010011;  // xori x12, x6, 12

        // // Shift immediate (I-type)
        // rom[26] = 32'b0000000_00101_00110_001_01101_0010011;  // slli x13, x6, 5
        // rom[27] = 32'b0000000_00001_00110_101_01110_0010011;  // srli x14, x6, 1
        // rom[28] = 32'b0100000_00010_00110_101_01111_0010011;  // srai x15, x6, 2

        // // U-type            
        // rom[29] = 32'b00000000000000000001_00101_0110111;  // LUI   x5, 0x1
        // rom[30] = 32'b00000000000000000010_00110_0010111;  // AUIPC x6, 0x2

        // // J-type
        // // rd = PC+4; PC += imm
        // rom[31] = 32'b000000000001_00000000_0000_00001_1101111;  // JAL  x16, 16
        
        // // rd = PC+4; PC = rs1 + imm
         rom[35] = 32'b00000000100000000000001001100111;      // JALR x4, 8(x0)    8+x0 = 8 -> 8/4  = 2번지로
        
    end



    assign inst_code = rom[inst_read_addr[31:2]];

endmodule
